`define RNOP    3'b111
`define RADD    3'b000
`define RSUB    3'b001
`define RMUL    3'b010
`define RB      3'b011
//`define ROR     3'b100
//`define RXOR    3'b101
//`define RNOR    3'b110